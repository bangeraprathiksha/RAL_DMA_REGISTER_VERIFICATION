`define no_of_trans 5


package ral_pkg;

  import uvm_pkg::*;
  `include "uvm_macros.svh"

	`include "defines.sv"

  // registers
  `include "registers.sv"

  // register block
  `include "top_reg_block.sv"

   // sequence item
  `include "reg_seq_item.sv"

  // sequence
  `include "top_reg_seq.sv"

  // driver
  `include "driver.sv"

  // monitor
  `include "monitor.sv"

  // adapter
  `include "adapter.sv"

  //agent
  `include "agent.sv"

  // environment
  `include "env.sv"

  // test
  `include "test.sv"

endpackage
